module display_module();
endmodule