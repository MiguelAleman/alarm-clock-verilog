module datapath(output [6:0] hours1, hours0, mins1, mins0, days, output am, pm, dblink, sound, input Next, Up, Set_Time, Set_Alarm, Snooze, Stop, Mute, Reset, Clr, Clk);
	// Control Units
		
endmodule